`timescale 1ns/10ps

module PriorityEncoder (P2, P1, P0, I7, I6, I5, I4, I3, I2, I1, I0);
	input I0, I1, I2, I3, I4, I5, I6, I7;
	output P2, P1, P0;
	wire I7I6, I6I5, I5I4, I6I5B, I6I5BI4, I6I5I4, I3I2; 
	wire I7B, I5B, I7I6B, I7BI7I6BI5B, I3B, I2B, I2BI1, I6I5I4I3BI2BI1, P0B;
	
	//P2
	NOR2X1 nor1(I7I6, I7, I6); //also used for P1 & P0
	NOR2X1 nor2(I5I4, I5, I4);
	NAND2X1 nand1(P2, I7I6, I5I4);
	
	//P1
	NOR2X1 nor3(I6I5, I6, I5);
	INVX2 inv1(I6I5B, I6I5);
	NOR2X1 nor4(I6I5BI4, I6I5B, I4);
	INVX2 inv2 (I6I5I4, I6I5BI4); //also used for P0
	NOR2X1 nor5(I3I2, I3, I2);
	OAI21X1 oai1(P1, I7I6, I6I5I4, I3I2);
	
	//P0
	INVX2 inv3(I7B, I7);
	INVX2 inv4(I5B, I5);
	INVX2 inv5(I7I6B, I7I6);
	OAI21X1 oai2(I7BI7I6BI5B, I7B, I7I6B, I5B);
	INVX2 inv6(I3B, I3);
	INVX2 inv7(I2B, I2);
	NAND2X1 nand2(I2BI1, I2B, I1);
	AOI21X1 aoi1(I6I5I4I3BI2BI1, I6I5I4, I3B, I2BI1);
	NOR2X1 nor6(P0B, I7BI7I6BI5B, I6I5I4I3BI2BI1);
	INVX2 inv8(P0, P0B);
endmodule