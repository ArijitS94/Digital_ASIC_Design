module AND2X1 (y, a, b);
	input a, b;
	output y;
	assign y = a & b;
endmodule

module OR2X1 (y, a, b);
	input a, b;
	output y;
	assign y = a | b;
endmodule

